module apple_tb();
	
	
	
endmodule
